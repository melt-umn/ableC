grammar edu:umn:cs:melt:exts:ableC:matrix;

exports edu:umn:cs:melt:exts:ableC:matrix:matrixSyntax;
exports edu:umn:cs:melt:exts:ableC:matrix:matrixStmt;
exports edu:umn:cs:melt:exts:ableC:matrix:matrixExpr;

