grammar edu:umn:cs:melt:ableC:abstractsyntax;

imports silver:langutil;
imports silver:langutil:pp;
imports edu:umn:cs:melt:ableC:abstractsyntax:env;
imports edu:umn:cs:melt:ableC:abstractsyntax:construction;

-- This module adds a new synthesized attribute that does not depend on the forward,
-- so it must be exported.  
exports edu:umn:cs:melt:ableC:abstractsyntax:substitution;
