grammar edu:umn:cs:melt:exts:ableC:adt;

exports edu:umn:cs:melt:exts:ableC:adt:concretesyntax:datatype;
exports edu:umn:cs:melt:exts:ableC:adt:concretesyntax:datatypeFwd;
exports edu:umn:cs:melt:exts:ableC:adt:concretesyntax:matchConstruct;
exports edu:umn:cs:melt:exts:ableC:adt:concretesyntax:matchConstructExpr;

exports edu:umn:cs:melt:exts:ableC:adt:abstractsyntax;
