grammar edu:umn:cs:melt:exts:ableC:closure;

exports edu:umn:cs:melt:exts:ableC:closure:concretesyntax:lambdaExpr;
exports edu:umn:cs:melt:exts:ableC:closure:concretesyntax:typeExpr;

exports edu:umn:cs:melt:exts:ableC:closure:abstractsyntax;