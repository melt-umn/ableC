grammar edu:umn:cs:melt:ableC:silverconstruction;

exports edu:umn:cs:melt:ableC:silverconstruction:concretesyntax;
