grammar edu:umn:cs:melt:exts:ableC:tables;

exports edu:umn:cs:melt:exts:ableC:tables:tableExpr;

