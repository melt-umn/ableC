grammar artifact;

import edu:umn:cs:melt:ableC:drivers:compile;

-- TODO: MDA test for this artifact

construct ableC as
edu:umn:cs:melt:ableC:concretesyntax
translator using
  edu:umn:cs:melt:tutorials:ableC:tainted;

