grammar edu:umn:cs:melt:exts:ableC:string:mda_test;

import edu:umn:cs:melt:ableC:host;

copper_mda testLambdaExpr(ablecParser) {
  edu:umn:cs:melt:exts:ableC:string:concretesyntax:str;
}

copper_mda testLambdaExpr(ablecParser) {
  edu:umn:cs:melt:exts:ableC:string:concretesyntax:show;
}

copper_mda testLambdaExpr(ablecParser) {
  edu:umn:cs:melt:exts:ableC:string:concretesyntax:typeExpr;
}