grammar edu:umn:cs:melt:exts:ableC:regex;

-- To make it as easy as including :regex into the parser, we export each bit of syntax from this grammar.
exports edu:umn:cs:melt:exts:ableC:regex:regexLiterals;
exports edu:umn:cs:melt:exts:ableC:regex:regexMatching;

