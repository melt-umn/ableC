
aspect production eqExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}
aspect production mulEqExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}
aspect production divEqExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}
aspect production modEqExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}
aspect production addEqExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}
aspect production subEqExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}
aspect production lshEqExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}
aspect production rshEqExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}
aspect production andEqExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}
aspect production orEqExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}
aspect production xorEqExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}



aspect production andExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}
aspect production orExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}



aspect production andBitExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}
aspect production orBitExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}
aspect production xorExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}
aspect production lshExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}
aspect production rshExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}



aspect production equalsExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}
aspect production notEqualsExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}
aspect production gtExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}
aspect production ltExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}
aspect production gteExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}
aspect production lteExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}

aspect production addExpr
top::Expr ::= lhs::Expr  rhs::Expr
{
  propagate substituted;
}
aspect production subExpr
top::Expr ::= lhs::Expr  rhs::Expr
{
  propagate substituted;
}
aspect production mulExpr
top::Expr ::= lhs::Expr  rhs::Expr
{
  propagate substituted;
}
aspect production divExpr
top::Expr ::= lhs::Expr  rhs::Expr
{
  propagate substituted;
}
aspect production modExpr
top::Expr ::= lhs::Expr  rhs::Expr
{
  propagate substituted;
}

aspect production commaExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}


aspect production ovrld:eqExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}
aspect production ovrld:mulEqExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}
aspect production ovrld:divEqExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}
aspect production ovrld:modEqExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}
aspect production ovrld:addEqExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}
aspect production ovrld:subEqExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}
aspect production ovrld:lshEqExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}
aspect production ovrld:rshEqExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}
aspect production ovrld:andEqExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}
aspect production ovrld:orEqExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}
aspect production ovrld:xorEqExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}



aspect production ovrld:andExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}
aspect production ovrld:orExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}



aspect production ovrld:andBitExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}
aspect production ovrld:orBitExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}
aspect production ovrld:xorExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}
aspect production ovrld:lshExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}
aspect production ovrld:rshExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}



aspect production ovrld:equalsExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}
aspect production ovrld:notEqualsExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}
aspect production ovrld:gtExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}
aspect production ovrld:ltExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}
aspect production ovrld:gteExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}
aspect production ovrld:lteExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}

aspect production ovrld:addExpr
top::Expr ::= lhs::Expr  rhs::Expr
{
  propagate substituted;
}
aspect production ovrld:subExpr
top::Expr ::= lhs::Expr  rhs::Expr
{
  propagate substituted;
}
aspect production ovrld:mulExpr
top::Expr ::= lhs::Expr  rhs::Expr
{
  propagate substituted;
}
aspect production ovrld:divExpr
top::Expr ::= lhs::Expr  rhs::Expr
{
  propagate substituted;
}
aspect production ovrld:modExpr
top::Expr ::= lhs::Expr  rhs::Expr
{
  propagate substituted;
}


aspect production inj:eqExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}
aspect production inj:mulEqExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}
aspect production inj:divEqExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}
aspect production inj:modEqExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}
aspect production inj:addEqExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}
aspect production inj:subEqExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}
aspect production inj:lshEqExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}
aspect production inj:rshEqExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}
aspect production inj:andEqExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}
aspect production inj:orEqExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}
aspect production inj:xorEqExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}



aspect production inj:andExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}
aspect production inj:orExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}



aspect production inj:andBitExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}
aspect production inj:orBitExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}
aspect production inj:xorExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}
aspect production inj:lshExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}
aspect production inj:rshExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}



aspect production inj:equalsExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}
aspect production inj:notEqualsExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}
aspect production inj:gtExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}
aspect production inj:ltExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}
aspect production inj:gteExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}
aspect production inj:lteExpr
top::Expr ::= lhs::Expr rhs::Expr
{
  propagate substituted;
}

aspect production inj:addExpr
top::Expr ::= lhs::Expr  rhs::Expr
{
  propagate substituted;
}
aspect production inj:subExpr
top::Expr ::= lhs::Expr  rhs::Expr
{
  propagate substituted;
}
aspect production inj:mulExpr
top::Expr ::= lhs::Expr  rhs::Expr
{
  propagate substituted;
}
aspect production inj:divExpr
top::Expr ::= lhs::Expr  rhs::Expr
{
  propagate substituted;
}
aspect production inj:modExpr
top::Expr ::= lhs::Expr  rhs::Expr
{
  propagate substituted;
}

