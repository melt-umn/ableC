grammar edu:umn:cs:melt:tutorials:ableC:helloworld;

exports edu:umn:cs:melt:tutorials:ableC:helloworld:abstractsyntax;
exports edu:umn:cs:melt:tutorials:ableC:helloworld:concretesyntax;