
synthesized attribute maybeRefId::Maybe<String> occurs on Attributes, Attribute, Attribs, Attrib;
attribute moduleName occurs on Attributes, Attribute, Attribs, Attrib;

synthesized attribute isHostAttrib::Boolean occurs on Attrib;

