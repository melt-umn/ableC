
fun fromId Name ::= n::cst:Identifier_t = name(n.lexeme);
fun fromTy Name ::= n::cst:TypeName_t = name(n.lexeme);

