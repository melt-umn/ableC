grammar edu:umn:cs:melt:exts:ableC:vector:mda_test;

import edu:umn:cs:melt:ableC:host;

--copper_mda testLambdaExpr(ablecParser) {
--  edu:umn:cs:melt:exts:ableC:vector:concretesyntax:constructor;
--}

copper_mda testLambdaExpr(ablecParser) {
  edu:umn:cs:melt:exts:ableC:vector:concretesyntax:typeExpr;
}