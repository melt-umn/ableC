grammar edu:umn:cs:melt:ableC:silverconstruction:concretesyntax;

exports edu:umn:cs:melt:ableC:silverconstruction:concretesyntax:quotation;
exports edu:umn:cs:melt:ableC:silverconstruction:concretesyntax:antiquotation;

exports edu:umn:cs:melt:ableC:concretesyntax;
exports edu:umn:cs:melt:ableC:concretesyntax:construction;
