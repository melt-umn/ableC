grammar edu:umn:cs:melt:exts:ableC:vector:mda_test;

import edu:umn:cs:melt:ableC:host;

--copper_mda testConstructor(ablecParser) {
--  edu:umn:cs:melt:exts:ableC:vector:concretesyntax:constructor;
--}

copper_mda testTypeExpr(ablecParser) {
  edu:umn:cs:melt:exts:ableC:vector:concretesyntax:typeExpr;
}