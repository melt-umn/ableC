grammar edu:umn:cs:melt:exts:ableC:adt:concretesyntax:matchKeyword;

imports edu:umn:cs:melt:ableC:concretesyntax;

marking terminal Match_t 'match' lexer classes {Ckeyword};


