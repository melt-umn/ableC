grammar edu:umn:cs:melt:ableC:host;

imports edu:umn:cs:melt:ableC:concretesyntax as cst;

parser ablecParser :: cst:Root {
  edu:umn:cs:melt:ableC:concretesyntax;
}

