grammar edu:umn:cs:melt:tutorials:ableC:tainted;

exports edu:umn:cs:melt:tutorials:ableC:tainted:abstractsyntax;
exports edu:umn:cs:melt:tutorials:ableC:tainted:concretesyntax;
