grammar edu:umn:cs:melt:ableC:abstractsyntax;

imports silver:langutil;
imports silver:langutil:pp;
imports edu:umn:cs:melt:ableC:abstractsyntax:env;
imports edu:umn:cs:melt:ableC:abstractsyntax:construction;

option edu:umn:cs:melt:ableC:abstractsyntax:substitution; -- TODO: Should this be an export?
