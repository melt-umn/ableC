grammar edu:umn:cs:melt:exts:ableC:templating;

exports edu:umn:cs:melt:exts:ableC:templating:concretesyntax;
exports edu:umn:cs:melt:exts:ableC:templating:abstractsyntax;