grammar edu:umn:cs:melt:exts:ableC:templating:mda_test;

import edu:umn:cs:melt:ableC:host;
{- TODO: FIX
copper_mda testTemplateDecl(ablecParser) {
  edu:umn:cs:melt:exts:ableC:templating:concretesyntax:templateDecl;
}

copper_mda testUsingDecl(ablecParser) {
  edu:umn:cs:melt:exts:ableC:templating:concretesyntax:templateDecl;
}
-}

copper_mda testInstExpr(ablecParser) {
  edu:umn:cs:melt:exts:ableC:templating:concretesyntax:instantiationExpr;
}

copper_mda testInstTypeExpr(ablecParser) {
  edu:umn:cs:melt:exts:ableC:templating:concretesyntax:instantiationTypeExpr;
}