grammar edu:umn:cs:melt:exts:ableC:gc;

-- To make it as easy as including :gc into the parser, we export each bit of syntax from this grammar.
exports edu:umn:cs:melt:exts:ableC:gc:gcMalloc;
exports edu:umn:cs:melt:exts:ableC:gc:gcRealloc;
exports edu:umn:cs:melt:exts:ableC:gc:gcNew;
