grammar edu:umn:cs:melt:exts:ableC:string;

exports edu:umn:cs:melt:exts:ableC:string:concretesyntax:typeExpr;
exports edu:umn:cs:melt:exts:ableC:string:concretesyntax:constructor;
exports edu:umn:cs:melt:exts:ableC:string:abstractsyntax;