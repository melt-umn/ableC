grammar edu:umn:cs:melt:exts:ableC:templating:mda_test;

import edu:umn:cs:melt:ableC:host;

copper_mda testDecl(ablecParser) {
  edu:umn:cs:melt:exts:ableC:templating:concretesyntax:templateDecl;
}

copper_mda testInstExpr(ablecParser) {
  edu:umn:cs:melt:exts:ableC:templating:concretesyntax:instantiationExpr;
}

copper_mda testInstTypeExpr(ablecParser) {
  edu:umn:cs:melt:exts:ableC:templating:concretesyntax:instantiationTypeExpr;
}