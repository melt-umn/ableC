grammar edu:umn:cs:melt:exts:silver:ableC:mda_test;

import silver:composed:Default;

copper_mda testAbleCEmbed(svParse) {
  edu:umn:cs:melt:exts:silver:ableC:concretesyntax;
}
