
abstract production extensionGenerated
top::OriginNote ::= string::String
{
  
}