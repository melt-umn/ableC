grammar edu:umn:cs:melt:exts:ableC:string;

exports edu:umn:cs:melt:exts:ableC:string:concretesyntax:typeExpr;
exports edu:umn:cs:melt:exts:ableC:string:concretesyntax:show;
exports edu:umn:cs:melt:exts:ableC:string:abstractsyntax;