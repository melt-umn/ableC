grammar edu:umn:cs:melt:exts:ableC:mex;

-- To make it as easy as including :mex into the parser, we export each bit of syntax from this grammar.
exports edu:umn:cs:melt:exts:ableC:mex:mexfunction;

-- We also depend upon the matrix extension's 'matrix' indexing syntax
exports edu:umn:cs:melt:exts:ableC:matrix:matrixSyntax;
exports edu:umn:cs:melt:exts:ableC:matrix:matrixExpr;

