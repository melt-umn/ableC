grammar edu:umn:cs:melt:tutorials:ableC:exponent;

exports edu:umn:cs:melt:tutorials:ableC:exponent:abstractsyntax;
exports edu:umn:cs:melt:tutorials:ableC:exponent:concretesyntax;