grammar edu:umn:cs:melt:exts:ableC:parfor;

exports edu:umn:cs:melt:exts:ableC:parfor:concretesyntax;

