grammar edu:umn:cs:melt:tutorials:ableC:globalint;

exports edu:umn:cs:melt:tutorials:ableC:globalint:abstractsyntax;
exports edu:umn:cs:melt:tutorials:ableC:globalint:concretesyntax;