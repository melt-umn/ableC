grammar edu:umn:cs:melt:exts:ableC:closure;

imports edu:umn:cs:melt:exts:ableC:gc;

exports edu:umn:cs:melt:exts:ableC:closure:concretesyntax:lambdaExpr;
exports edu:umn:cs:melt:exts:ableC:closure:concretesyntax:typeExpr;

exports edu:umn:cs:melt:exts:ableC:closure:abstractsyntax;