grammar edu:umn:cs:melt:exts:ableC:adt:mda_test;

import edu:umn:cs:melt:ableC:host;

copper_mda testDatatype(ablecParser) {
  edu:umn:cs:melt:exts:ableC:gcadt:concretesyntax:datatype;
}