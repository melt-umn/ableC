grammar edu:umn:cs:melt:tutorials:ableC:tuple;

exports edu:umn:cs:melt:tutorials:ableC:tuple:abstractsyntax;
exports edu:umn:cs:melt:tutorials:ableC:tuple:concretesyntax;