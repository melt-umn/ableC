grammar edu:umn:cs:melt:tutorials:ableC:average;

exports edu:umn:cs:melt:tutorials:ableC:average:abstractsyntax;
exports edu:umn:cs:melt:tutorials:ableC:average:concretesyntax;