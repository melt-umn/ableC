grammar edu:umn:cs:melt:exts:ableC:vector;

exports edu:umn:cs:melt:exts:ableC:vector:concretesyntax:typeExpr;
exports edu:umn:cs:melt:exts:ableC:vector:concretesyntax:constructor;

exports edu:umn:cs:melt:exts:ableC:vector:abstractsyntax;