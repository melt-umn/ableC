grammar edu:umn:cs:melt:tutorials:ableC:interval:concretesyntax;

exports edu:umn:cs:melt:tutorials:ableC:interval:concretesyntax:typeExpr;
exports edu:umn:cs:melt:tutorials:ableC:interval:concretesyntax:constructor;