grammar edu:umn:cs:melt:exts:ableC:matrix:mda_test;

import edu:umn:cs:melt:ableC:host;

copper_mda testStmt(ablecParser) {
  edu:umn:cs:melt:exts:ableC:matrix:matrixSyntax;
  edu:umn:cs:melt:exts:ableC:matrix:matrixStmt;
}

copper_mda testExpr(ablecParser) {
  edu:umn:cs:melt:exts:ableC:matrix:matrixSyntax;
  edu:umn:cs:melt:exts:ableC:matrix:matrixExpr;
}

