grammar edu:umn:cs:melt:exts:ableC:regex;

import edu:umn:cs:melt:ableC:host;

copper_mda testMatching(ablecParser) {
  edu:umn:cs:melt:exts:ableC:regex:regexMatching;
}

copper_mda testLiterals(ablecParser) {
  edu:umn:cs:melt:exts:ableC:regex:regexLiterals;
}

