grammar edu:umn:cs:melt:tutorials:ableC:intconst;

exports edu:umn:cs:melt:tutorials:ableC:intconst:abstractsyntax;
exports edu:umn:cs:melt:tutorials:ableC:intconst:concretesyntax;