grammar edu:umn:cs:melt:exts:ableC:tables:mda_test;

import edu:umn:cs:melt:ableC:host;

copper_mda testTables(ablecParser) {
  edu:umn:cs:melt:exts:ableC:tables:tableExpr;
}

