grammar edu:umn:cs:melt:tutorials:ableC:interval;

exports edu:umn:cs:melt:tutorials:ableC:interval:abstractsyntax;
exports edu:umn:cs:melt:tutorials:ableC:interval:concretesyntax;