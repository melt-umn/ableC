grammar edu:umn:cs:melt:exts:ableC:adt:mda_test;

import edu:umn:cs:melt:ableC:host;

copper_mda testMatchStmt(ablecParser) {
  edu:umn:cs:melt:exts:ableC:adt:concretesyntax:matchConstruct;
}
copper_mda testMatchExpr(ablecParser) {
  edu:umn:cs:melt:exts:ableC:adt:concretesyntax:matchConstructExpr;
}
copper_mda testDatatype(ablecParser) {
  edu:umn:cs:melt:exts:ableC:adt:concretesyntax:datatype;
}
copper_mda testDatatypeFwd(ablecParser) {
  edu:umn:cs:melt:exts:ableC:adt:concretesyntax:datatypeFwd;
}

