grammar edu:umn:cs:melt:ableC:abstractsyntax:substitution;


synthesized attribute host<a>::a;