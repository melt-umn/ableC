grammar edu:umn:cs:melt:ableC:abstractsyntax;

synthesized attribute host<a>::a;