grammar edu:umn:cs:melt:tutorials:ableC:prefixExpr;

exports edu:umn:cs:melt:tutorials:ableC:prefixExpr:abstractsyntax;
exports edu:umn:cs:melt:tutorials:ableC:prefixExpr:concretesyntax;