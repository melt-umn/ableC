grammar edu:umn:cs:melt:ableC:abstractsyntax;

imports silver:langutil;
imports silver:langutil:pp with implode as ppImplode;
imports edu:umn:cs:melt:ableC:abstractsyntax:env;

