grammar edu:umn:cs:melt:exts:ableC:mex:mda_test;

import edu:umn:cs:melt:ableC:host;

copper_mda testMex(ablecParser) {
  edu:umn:cs:melt:exts:ableC:mex:mexfunction;
}


