grammar edu:umn:cs:melt:exts:ableC:closure:mda_test;

import edu:umn:cs:melt:ableC:host;

copper_mda testLambdaExpr(ablecParser) {
  edu:umn:cs:melt:exts:ableC:closure:concretesyntax:lambdaExpr;
}

copper_mda testTypeExpr(ablecParser) {
  edu:umn:cs:melt:exts:ableC:closure:concretesyntax:typeExpr;
}

