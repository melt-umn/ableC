grammar edu:umn:cs:melt:exts:silver:ableC;

exports edu:umn:cs:melt:exts:silver:ableC:concretesyntax;
